module hk(output ed);
  assign ed=1;
endmodule
