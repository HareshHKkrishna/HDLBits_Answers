module test
  test to streak;
endmodule
